module axi_crossbar_wr #
(
    parameter M_REGIONS= 1,
    parameter S_IF_COUNT = 4,
    parameter M_IF_COUNT = 4,
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 32,
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    parameter S_IF_ID_WIDTH = 8,
    parameter M_IF_ID_WIDTH = S_IF_ID_WIDTH+$clog2(S_IF_COUNT),
    parameter M_BASE_ADDR = 0,
    parameter M_ADDR_WIDTH = {M_IF_COUNT{{M_REGIONS{32'd24}}}},
    parameter M_CONNECT = {M_IF_COUNT{{S_IF_COUNT{1'b1}}}},
    parameter S_AW_FIFO = {S_IF_COUNT{2'd0}},
    parameter S_W_FIFO = {S_IF_COUNT{2'd0}},
    parameter S_B_FIFO = {S_IF_COUNT{2'd1}},
    parameter M_AW_FIFO = {M_IF_COUNT{2'd1}},
    parameter M_W_FIFO = {M_IF_COUNT{2'd2}},
    parameter M_B_FIFO = {M_IF_COUNT{2'd0}}
)
(
    input                                 clk,
    input                                 rst,
    input  [S_IF_COUNT*S_IF_ID_WIDTH-1:0] s_axi_awid,
    input  [S_IF_COUNT*ADDR_WIDTH-1:0]    s_axi_awaddr,
    input  [S_IF_COUNT*8-1:0]             s_axi_awlen,
    input  [S_IF_COUNT*3-1:0]             s_axi_awsize,
    input  [S_IF_COUNT*2-1:0]             s_axi_awburst,
    input  [S_IF_COUNT-1:0]               s_axi_awlock,
    input  [S_IF_COUNT*4-1:0]             s_axi_awqos,
    input  [S_IF_COUNT-1:0]               s_axi_awvalid,
    output [S_IF_COUNT-1:0]               s_axi_awready,
    input  [S_IF_COUNT*S_IF_ID_WIDTH-1:0] s_axi_wid,
    input  [S_IF_COUNT*DATA_WIDTH-1:0]    s_axi_wdata,
    input  [S_IF_COUNT*STRB_WIDTH-1:0]    s_axi_wstrb,
    input  [S_IF_COUNT-1:0]               s_axi_wlast,
    input  [S_IF_COUNT-1:0]               s_axi_wvalid,
    output [S_IF_COUNT-1:0]               s_axi_wready,
    output [S_IF_COUNT*S_IF_ID_WIDTH-1:0] s_axi_bid,
    output [S_IF_COUNT*2-1:0]             s_axi_bresp,
    output [S_IF_COUNT-1:0]               s_axi_bvalid,
    input  [S_IF_COUNT-1:0]               s_axi_bready,
    output [M_IF_COUNT*M_IF_ID_WIDTH-1:0] m_axi_awid,
    output [M_IF_COUNT*ADDR_WIDTH-1:0]    m_axi_awaddr,
    output [M_IF_COUNT*8-1:0]             m_axi_awlen,
    output [M_IF_COUNT*3-1:0]             m_axi_awsize,
    output [M_IF_COUNT*2-1:0]             m_axi_awburst,
    output [M_IF_COUNT-1:0]               m_axi_awlock,
    output [M_IF_COUNT*4-1:0]             m_axi_awqos,
    output [M_IF_COUNT-1:0]               m_axi_awvalid,
    input  [M_IF_COUNT-1:0]               m_axi_awready,
    output [M_IF_COUNT*M_IF_ID_WIDTH-1:0] m_axi_wid,
    output [M_IF_COUNT*DATA_WIDTH-1:0]    m_axi_wdata,
    output [M_IF_COUNT*STRB_WIDTH-1:0]    m_axi_wstrb,
    output [M_IF_COUNT-1:0]               m_axi_wlast,
    output [M_IF_COUNT-1:0]               m_axi_wvalid,
    input  [M_IF_COUNT-1:0]               m_axi_wready,
    input  [M_IF_COUNT*M_IF_ID_WIDTH-1:0] m_axi_bid,
    input  [M_IF_COUNT*2-1:0]             m_axi_bresp,
    input  [M_IF_COUNT-1:0]               m_axi_bvalid,
    output [M_IF_COUNT-1:0]               m_axi_bready,

    output [S_IF_COUNT*ADDR_WIDTH-1:0]    wr_error_addr,
    output [S_IF_COUNT-1:0]               wr_error_valid,
    input  [S_IF_COUNT-1:0]               wr_error_ready
);
endmodule