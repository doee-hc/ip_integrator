`define  ARBITER_WIDTH 3
`define  PORTS `ARBITER_WIDTH
