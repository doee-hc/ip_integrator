`include "arbiter_config_0.vh"

`define  ARBITER_WIDTH 5
`define  PORTS `ARBITER_WIDTH

`define  ARB_BLOCK_ACK 1

`define  ARB_LSB_HIGH_PRIORITY
