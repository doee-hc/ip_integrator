

`timescale 1ns / 1ps

//------------------------------------------------------------------------------
// Module
//------------------------------------------------------------------------------

module litespi_core_axi_lite (
    input  wire   [31:0] bus_araddr,
    input  wire    [2:0] bus_arprot,
    output wire          bus_arready,
    input  wire          bus_arvalid,
    input  wire   [31:0] bus_awaddr,
    input  wire    [2:0] bus_awprot,
    output wire          bus_awready,
    input  wire          bus_awvalid,
    input  wire          bus_bready,
    output wire    [1:0] bus_bresp,
    output wire          bus_bvalid,
    output wire   [31:0] bus_rdata,
    input  wire          bus_rready,
    output wire    [1:0] bus_rresp,
    output wire          bus_rvalid,
    input  wire   [31:0] bus_wdata,
    output wire          bus_wready,
    input  wire    [3:0] bus_wstrb,
    input  wire          bus_wvalid,
    input  wire          clk,
    input  wire          rst,
    output reg           spiflash_clk,
    output wire          spiflash_cs_n,
    input  wire          spiflash_hold,
    input  wire          spiflash_miso,
    output reg           spiflash_mosi,
    input  wire          spiflash_wp
);



//------------------------------------------------------------------------------
// Specialized Logic
//------------------------------------------------------------------------------

endmodule

// -----------------------------------------------------------------------------
//  Auto-Generated by LiteX on 2024-06-15 18:04:14.
//------------------------------------------------------------------------------
