`define  ARBITER_WIDTH 4
`define  PORTS `ARBITER_WIDTH
